module debouncer (

);

endmodule