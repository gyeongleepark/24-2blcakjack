`timescale 1ns / 1ps

module top(
    input clk,
    input reset,
    input next,
    input hit,
    input stand,
    input double,
    input split,
    input bet_8,
    input bet_4,
    input bet_2,
    input bet_1,
    output reg [5:0] player_current_score,      // Final player score
    output reg [5:0] player_new_card,          // Latest player card
    output reg [5:0] player_current_score_split, // Score for split hand
    output reg [5:0] player_new_card_split,    // Latest split hand card
    output reg [5:0] dealer_current_score,     // Final dealer score
    output reg [4:0] current_coin,             // Player's current coins
    output reg can_split,                      // Indicates if split is possible
    output reg Win,                            // Win flag
    output reg Lose,                           // Lose flag
    output reg Draw                            // Draw flag
);

    // Internal signals
    reg [2:0] game_state;                   // Tracks the game phase (e.g., betting, dealing, result)
    reg [5:0] player_hand [1:4];            // Player's cards (up to 4 cards per hand)
    reg [5:0] dealer_hand [1:4];            // Dealer's cards (up to 4 cards)
    reg [5:0] split_hand [1:4];             // Player's split hand cards
    reg [1:0] hand_count;                   // Number of player hands (used for splits)
    reg [3:0] player_card_count, dealer_card_count, split_card_count; // Card counts for each hand

    reg [5:0] player_score_internal;        // Internal score for player's main hand
    reg [5:0] dealer_score_internal;        // Internal score for dealer
    reg [5:0] split_score_internal;         // Internal score for split hand
    reg [4:0] coin_internal;                // Internal coin count
    reg split_flag_internal;                // Indicates if split was activated
    reg win_flag_internal, lose_flag_internal, draw_flag_internal; // Result flags

    wire [3:0] card1, card2;                // Cards generated by card_generation module

    // Card generation module instantiation
    card_generation card_gen (
        .clk(clk),
        .reset(reset),
        .on(next),                          // Generate new cards on "next"
        .test(3'b000),                      // Change to desired test case
        .card1_out(card1),
        .card2_out(card2)
    );

    // Game states
    localparam STATE_BETTING    = 3'b000,
               STATE_DEALER_CARD = 3'b001,
               STATE_PLAYER_CARD = 3'b010,
               STATE_SPLIT       = 3'b011,
               STATE_RESULT      = 3'b100;

    // Clock-driven behavior
    always @(posedge clk or posedge reset) begin
        if (reset) begin
            // Initialize all signals
            game_state <= STATE_BETTING;
            player_card_count <= 0;
            dealer_card_count <= 0;
            split_card_count <= 0;
            hand_count <= 1;
            player_score_internal <= 0;
            dealer_score_internal <= 0;
            split_score_internal <= 0;
            coin_internal <= 5'd30;         // Start with 30 coins
            split_flag_internal <= 0;
            win_flag_internal <= 0;
            lose_flag_internal <= 0;
            draw_flag_internal <= 0;
        end else begin
            case (game_state)
                // Betting phase
                STATE_BETTING: begin
                    if (bet_8 || bet_4 || bet_2 || bet_1) begin      // 잔액 부족할 때 아직 모름
                        // Calculate bet amount and move to the next phase
                        // 총 베팅 금액 계산
                        reg [4:0] total_bet; // 총 베팅 금액 임시 저장 변수
                        total_bet = bet_8 * 8 + bet_4 * 4 + bet_2 * 2 + bet_1 * 1;

                        if (total_bet > 15) begin
                            // 베팅 금액이 최대 15를 초과하면, 15로 고정
                            coin_internal <= coin_internal - 15;
                        end else begin
                            // 그렇지 않으면 실제 베팅 금액 차감
                            coin_internal <= coin_internal - total_bet;
                        end

                        game_state <= STATE_DEALER_CARD;
                    end
                end

                // Dealer's initial card phase
                STATE_DEALER_CARD: begin
                    if (next) begin
                        dealer_hand[1] <= card1;
                        dealer_card_count <= 1;
                        dealer_score_internal <= card1;
                        game_state <= STATE_PLAYER_CARD;
                    end
                end

                // Player's initial card phase
                STATE_PLAYER_CARD: begin
                    if (next) begin
                        player_hand[1] <= card1;
                        player_hand[2] <= card2;
                        player_card_count <= 2;
                        player_score_internal <= card1 + card2;

                        // Check for split
                        if (card1 == card2)
                            split_flag_internal <= 1;

                        game_state <= STATE_SPLIT;
                    end
                end

                // Split handling phase
                STATE_SPLIT: begin
                    if (split && split_flag_internal) begin
                        hand_count <= 2; // Player now has two hands
                        split_hand[1] <= player_hand[2];
                        split_card_count <= 1;
                        player_card_count <= 1;
                        split_score_internal <= player_hand[2];
                        player_score_internal <= player_hand[1];
                    end else begin
                        game_state <= STATE_RESULT;
                    end
                end

                // Result phase
                STATE_RESULT: begin
                    if (player_score_internal > 21)
                        lose_flag_internal <= 1;
                    else if (dealer_score_internal > 21)
                        win_flag_internal <= 1;
                    else if (player_score_internal > dealer_score_internal)
                        win_flag_internal <= 1;
                    else if (player_score_internal < dealer_score_internal)
                        lose_flag_internal <= 1;
                    else
                        draw_flag_internal <= 1;
                end
            endcase
        end
    end

    // Output assignments
    always @(posedge clk or posedge reset) begin
        if (reset) begin
            player_current_score <= 0;
            dealer_current_score <= 0;
            player_new_card <= 0;
            player_current_score_split <= 0;
            player_new_card_split <= 0;
            current_coin <= 5'd10;
            can_split <= 0;
            Win <= 0;
            Lose <= 0;
            Draw <= 0;
        end else begin
            player_current_score <= player_score_internal;
            dealer_current_score <= dealer_score_internal;
            player_new_card <= player_hand[player_card_count];
            player_current_score_split <= split_score_internal;
            player_new_card_split <= split_hand[split_card_count];
            current_coin <= coin_internal;
            can_split <= split_flag_internal;
            Win <= win_flag_internal;
            Lose <= lose_flag_internal;
            Draw <= draw_flag_internal;
        end
    end

endmodule

/*
STATE_HIT: begin
    if (hit) begin
        // 카드 생성 모듈 활성화
        card_gen_enable <= 1;

        // 새로운 카드를 플레이어 핸드에 추가
        player_hand[player_card_count] <= card1;
        player_card_count <= player_card_count + 1;

        // 카드 생성 완료 후 모듈 비활성화
        card_gen_enable <= 0;

        // 버스트 여부 확인 (현재 점수가 21 초과)
        if ((player_current_score + card1) > 21) begin
            player_bust <= 1;
            game_state <= STATE_DEALER_TURN; // 딜러 턴으로 이동
        end
        else begin
            game_state <= STATE_HIT_STAND; // 플레이어가 추가로 hit/stand 선택
        end
    end
end

STATE_SPLIT: begin
    if (split && can_split) begin
        // 스플릿 처리
        split_active <= 1; // 스플릿 상태 활성화

        // 현재 첫 번째 카드만 남기고 분리
        player_split_hand[0] <= player_hand[1];
        player_card_count <= 1; // 현재 핸드는 첫 번째 카드만 유지

        // 두 번째 카드와 새 카드는 분리된 핸드로 처리
        player_hand_split[0] <= player_hand[2];
        player_hand_split[1] <= card1;
        split_card_count <= 2;

        // 다음 상태 설정
        game_state <= STATE_PLAYER_SPLIT; // 스플릿 핸드 처리 상태로 전이
    end
end

STATE_PLAYER_SPLIT: begin
    if (!split_done) begin
        if (hit_split) begin
            // 분리된 핸드에 추가 카드 지급
            player_hand_split[split_card_count] <= card1;
            split_card_count <= split_card_count + 1;

            // 버스트 여부 확인
            if ((player_current_score_split + card1) > 21) begin
                split_bust <= 1;
                game_state <= STATE_DEALER_TURN; // 딜러 턴으로 이동
            end
        end
        else if (stand_split) begin
            // 스탠드 선택 시 분리된 핸드 처리 완료
            split_done <= 1;
            game_state <= STATE_DEALER_TURN; // 딜러 턴으로 이동
        end
    end
end
*/